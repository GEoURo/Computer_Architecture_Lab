
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h610e9bbb;
    ram_cell[       1] = 32'h0;  // 32'hae80ab86;
    ram_cell[       2] = 32'h0;  // 32'h7ea90fdf;
    ram_cell[       3] = 32'h0;  // 32'h3a205879;
    ram_cell[       4] = 32'h0;  // 32'hf3190527;
    ram_cell[       5] = 32'h0;  // 32'hf706fd22;
    ram_cell[       6] = 32'h0;  // 32'hce019673;
    ram_cell[       7] = 32'h0;  // 32'h71a3c5bc;
    ram_cell[       8] = 32'h0;  // 32'h93cb1d7a;
    ram_cell[       9] = 32'h0;  // 32'h794fd1dc;
    ram_cell[      10] = 32'h0;  // 32'h84de14b8;
    ram_cell[      11] = 32'h0;  // 32'h7e1ae1b4;
    ram_cell[      12] = 32'h0;  // 32'h0ea2ddc2;
    ram_cell[      13] = 32'h0;  // 32'h219557a9;
    ram_cell[      14] = 32'h0;  // 32'hbb72d2c0;
    ram_cell[      15] = 32'h0;  // 32'h218867e3;
    ram_cell[      16] = 32'h0;  // 32'h8ccdee05;
    ram_cell[      17] = 32'h0;  // 32'hc5dc8973;
    ram_cell[      18] = 32'h0;  // 32'hdeabbeb6;
    ram_cell[      19] = 32'h0;  // 32'h7d8006f4;
    ram_cell[      20] = 32'h0;  // 32'h86d22415;
    ram_cell[      21] = 32'h0;  // 32'h5fdca60a;
    ram_cell[      22] = 32'h0;  // 32'h7ea4f82a;
    ram_cell[      23] = 32'h0;  // 32'h72a17ffc;
    ram_cell[      24] = 32'h0;  // 32'h33a0bc26;
    ram_cell[      25] = 32'h0;  // 32'h87948f58;
    ram_cell[      26] = 32'h0;  // 32'h29ded1c1;
    ram_cell[      27] = 32'h0;  // 32'h90959303;
    ram_cell[      28] = 32'h0;  // 32'h3d8ff206;
    ram_cell[      29] = 32'h0;  // 32'h5d25e7d2;
    ram_cell[      30] = 32'h0;  // 32'hc3b0125f;
    ram_cell[      31] = 32'h0;  // 32'hed95937d;
    ram_cell[      32] = 32'h0;  // 32'h18e6fac2;
    ram_cell[      33] = 32'h0;  // 32'h496b0f84;
    ram_cell[      34] = 32'h0;  // 32'heac99925;
    ram_cell[      35] = 32'h0;  // 32'h5fa7e47f;
    ram_cell[      36] = 32'h0;  // 32'h9b2cd279;
    ram_cell[      37] = 32'h0;  // 32'h329b1c8c;
    ram_cell[      38] = 32'h0;  // 32'hba94de49;
    ram_cell[      39] = 32'h0;  // 32'h2a83983c;
    ram_cell[      40] = 32'h0;  // 32'h5e28d4dc;
    ram_cell[      41] = 32'h0;  // 32'hea9d98b4;
    ram_cell[      42] = 32'h0;  // 32'hd0be81b8;
    ram_cell[      43] = 32'h0;  // 32'h22759e2e;
    ram_cell[      44] = 32'h0;  // 32'h0629516b;
    ram_cell[      45] = 32'h0;  // 32'h74606e7c;
    ram_cell[      46] = 32'h0;  // 32'h2b886838;
    ram_cell[      47] = 32'h0;  // 32'hb8614fbc;
    ram_cell[      48] = 32'h0;  // 32'h2262c3d2;
    ram_cell[      49] = 32'h0;  // 32'h9cbce6e4;
    ram_cell[      50] = 32'h0;  // 32'hfea44ff7;
    ram_cell[      51] = 32'h0;  // 32'h7ae3515a;
    ram_cell[      52] = 32'h0;  // 32'h13f98b73;
    ram_cell[      53] = 32'h0;  // 32'h9e2f63c3;
    ram_cell[      54] = 32'h0;  // 32'hdbc40723;
    ram_cell[      55] = 32'h0;  // 32'hd3dc5d15;
    ram_cell[      56] = 32'h0;  // 32'h76afe000;
    ram_cell[      57] = 32'h0;  // 32'h33503018;
    ram_cell[      58] = 32'h0;  // 32'hfa63496e;
    ram_cell[      59] = 32'h0;  // 32'h165f05c0;
    ram_cell[      60] = 32'h0;  // 32'h62fa3c23;
    ram_cell[      61] = 32'h0;  // 32'h21be49e9;
    ram_cell[      62] = 32'h0;  // 32'had54648c;
    ram_cell[      63] = 32'h0;  // 32'hb34572aa;
    ram_cell[      64] = 32'h0;  // 32'h999088cd;
    ram_cell[      65] = 32'h0;  // 32'h46c40ebb;
    ram_cell[      66] = 32'h0;  // 32'h21c46974;
    ram_cell[      67] = 32'h0;  // 32'h4ee4dd5c;
    ram_cell[      68] = 32'h0;  // 32'h4f9ec9b3;
    ram_cell[      69] = 32'h0;  // 32'h4db7aa83;
    ram_cell[      70] = 32'h0;  // 32'h66e4363b;
    ram_cell[      71] = 32'h0;  // 32'he56c6879;
    ram_cell[      72] = 32'h0;  // 32'hf53a5833;
    ram_cell[      73] = 32'h0;  // 32'hd43fc287;
    ram_cell[      74] = 32'h0;  // 32'hb0bd35d0;
    ram_cell[      75] = 32'h0;  // 32'h4a5dbc9c;
    ram_cell[      76] = 32'h0;  // 32'h0f5609b1;
    ram_cell[      77] = 32'h0;  // 32'hf250b301;
    ram_cell[      78] = 32'h0;  // 32'hedef4047;
    ram_cell[      79] = 32'h0;  // 32'ha4b77339;
    ram_cell[      80] = 32'h0;  // 32'hd34ae8d6;
    ram_cell[      81] = 32'h0;  // 32'h7ad102dd;
    ram_cell[      82] = 32'h0;  // 32'hfa212229;
    ram_cell[      83] = 32'h0;  // 32'h009ba3ce;
    ram_cell[      84] = 32'h0;  // 32'h25167bdd;
    ram_cell[      85] = 32'h0;  // 32'h5b10cda6;
    ram_cell[      86] = 32'h0;  // 32'hb1991060;
    ram_cell[      87] = 32'h0;  // 32'h2da67b55;
    ram_cell[      88] = 32'h0;  // 32'h413c2473;
    ram_cell[      89] = 32'h0;  // 32'hf7cde870;
    ram_cell[      90] = 32'h0;  // 32'h5971f742;
    ram_cell[      91] = 32'h0;  // 32'hdaf5c2ba;
    ram_cell[      92] = 32'h0;  // 32'hc9ab54d1;
    ram_cell[      93] = 32'h0;  // 32'h2bdb6f48;
    ram_cell[      94] = 32'h0;  // 32'h03187d8b;
    ram_cell[      95] = 32'h0;  // 32'hf0a81458;
    ram_cell[      96] = 32'h0;  // 32'h243561e3;
    ram_cell[      97] = 32'h0;  // 32'h7c77534c;
    ram_cell[      98] = 32'h0;  // 32'h26cff365;
    ram_cell[      99] = 32'h0;  // 32'h24712d79;
    ram_cell[     100] = 32'h0;  // 32'h54fe6d8e;
    ram_cell[     101] = 32'h0;  // 32'hb850955e;
    ram_cell[     102] = 32'h0;  // 32'ha413ac73;
    ram_cell[     103] = 32'h0;  // 32'h9f22361d;
    ram_cell[     104] = 32'h0;  // 32'h4b56a90f;
    ram_cell[     105] = 32'h0;  // 32'hb1105219;
    ram_cell[     106] = 32'h0;  // 32'hb6912cb0;
    ram_cell[     107] = 32'h0;  // 32'he71df1eb;
    ram_cell[     108] = 32'h0;  // 32'ha00e9a81;
    ram_cell[     109] = 32'h0;  // 32'h11f9220e;
    ram_cell[     110] = 32'h0;  // 32'h8e2c6132;
    ram_cell[     111] = 32'h0;  // 32'h7d46cb2e;
    ram_cell[     112] = 32'h0;  // 32'h15b6c243;
    ram_cell[     113] = 32'h0;  // 32'h4a36af0d;
    ram_cell[     114] = 32'h0;  // 32'hc1d0d442;
    ram_cell[     115] = 32'h0;  // 32'he6389145;
    ram_cell[     116] = 32'h0;  // 32'h85b5ffd3;
    ram_cell[     117] = 32'h0;  // 32'h480e6f92;
    ram_cell[     118] = 32'h0;  // 32'h82fc65b9;
    ram_cell[     119] = 32'h0;  // 32'hfb16c5a9;
    ram_cell[     120] = 32'h0;  // 32'h430bb8ec;
    ram_cell[     121] = 32'h0;  // 32'hdf7f2bb9;
    ram_cell[     122] = 32'h0;  // 32'hc36384d3;
    ram_cell[     123] = 32'h0;  // 32'h4ea71856;
    ram_cell[     124] = 32'h0;  // 32'h5fe309d2;
    ram_cell[     125] = 32'h0;  // 32'he0f940b3;
    ram_cell[     126] = 32'h0;  // 32'h87b16010;
    ram_cell[     127] = 32'h0;  // 32'hba797460;
    ram_cell[     128] = 32'h0;  // 32'h623bd4f3;
    ram_cell[     129] = 32'h0;  // 32'hb4753e52;
    ram_cell[     130] = 32'h0;  // 32'heb730f50;
    ram_cell[     131] = 32'h0;  // 32'h17c0201b;
    ram_cell[     132] = 32'h0;  // 32'h162dd68f;
    ram_cell[     133] = 32'h0;  // 32'h395d6a27;
    ram_cell[     134] = 32'h0;  // 32'h75205fa1;
    ram_cell[     135] = 32'h0;  // 32'hbb2b3619;
    ram_cell[     136] = 32'h0;  // 32'h1cc3ccc1;
    ram_cell[     137] = 32'h0;  // 32'hd08ad64b;
    ram_cell[     138] = 32'h0;  // 32'hb92b854e;
    ram_cell[     139] = 32'h0;  // 32'h203aaef5;
    ram_cell[     140] = 32'h0;  // 32'h56a3e721;
    ram_cell[     141] = 32'h0;  // 32'h7f54bd6b;
    ram_cell[     142] = 32'h0;  // 32'h918c9ba7;
    ram_cell[     143] = 32'h0;  // 32'h2b34bb32;
    ram_cell[     144] = 32'h0;  // 32'h1503c76e;
    ram_cell[     145] = 32'h0;  // 32'h02bd9f4f;
    ram_cell[     146] = 32'h0;  // 32'hd50faf43;
    ram_cell[     147] = 32'h0;  // 32'h8a3c4606;
    ram_cell[     148] = 32'h0;  // 32'h73005367;
    ram_cell[     149] = 32'h0;  // 32'h378e30ad;
    ram_cell[     150] = 32'h0;  // 32'hf0282dde;
    ram_cell[     151] = 32'h0;  // 32'h7cef0936;
    ram_cell[     152] = 32'h0;  // 32'hd1f1eb03;
    ram_cell[     153] = 32'h0;  // 32'hb41a9be8;
    ram_cell[     154] = 32'h0;  // 32'h3ad41b0f;
    ram_cell[     155] = 32'h0;  // 32'hf362e79e;
    ram_cell[     156] = 32'h0;  // 32'h15f27a98;
    ram_cell[     157] = 32'h0;  // 32'ha51b2d84;
    ram_cell[     158] = 32'h0;  // 32'ha1cb9673;
    ram_cell[     159] = 32'h0;  // 32'h0975cf13;
    ram_cell[     160] = 32'h0;  // 32'h8e17ce5d;
    ram_cell[     161] = 32'h0;  // 32'hf61d342b;
    ram_cell[     162] = 32'h0;  // 32'hbc787c7b;
    ram_cell[     163] = 32'h0;  // 32'h3d40c9d7;
    ram_cell[     164] = 32'h0;  // 32'h8e680a8a;
    ram_cell[     165] = 32'h0;  // 32'ha3ffdb29;
    ram_cell[     166] = 32'h0;  // 32'h43729b43;
    ram_cell[     167] = 32'h0;  // 32'h49a2e1a6;
    ram_cell[     168] = 32'h0;  // 32'hd52ce0ab;
    ram_cell[     169] = 32'h0;  // 32'h9ac441c6;
    ram_cell[     170] = 32'h0;  // 32'h671fd589;
    ram_cell[     171] = 32'h0;  // 32'hb5ae67cd;
    ram_cell[     172] = 32'h0;  // 32'he0410655;
    ram_cell[     173] = 32'h0;  // 32'h6b7a3341;
    ram_cell[     174] = 32'h0;  // 32'hee400bc3;
    ram_cell[     175] = 32'h0;  // 32'hc30b46ff;
    ram_cell[     176] = 32'h0;  // 32'h8acca5f9;
    ram_cell[     177] = 32'h0;  // 32'h94ec3172;
    ram_cell[     178] = 32'h0;  // 32'h85ba9a1c;
    ram_cell[     179] = 32'h0;  // 32'h79305390;
    ram_cell[     180] = 32'h0;  // 32'h90097457;
    ram_cell[     181] = 32'h0;  // 32'hb2b6ba33;
    ram_cell[     182] = 32'h0;  // 32'h5694fac1;
    ram_cell[     183] = 32'h0;  // 32'h98389cdc;
    ram_cell[     184] = 32'h0;  // 32'hcae7fe67;
    ram_cell[     185] = 32'h0;  // 32'h7ff0e0af;
    ram_cell[     186] = 32'h0;  // 32'hed8452e6;
    ram_cell[     187] = 32'h0;  // 32'h7c02aecb;
    ram_cell[     188] = 32'h0;  // 32'h07cac0af;
    ram_cell[     189] = 32'h0;  // 32'h6f9bd126;
    ram_cell[     190] = 32'h0;  // 32'hc3848f34;
    ram_cell[     191] = 32'h0;  // 32'h6e56618c;
    ram_cell[     192] = 32'h0;  // 32'h52404517;
    ram_cell[     193] = 32'h0;  // 32'h1676d525;
    ram_cell[     194] = 32'h0;  // 32'h40ad633d;
    ram_cell[     195] = 32'h0;  // 32'h01443334;
    ram_cell[     196] = 32'h0;  // 32'h1125961f;
    ram_cell[     197] = 32'h0;  // 32'he608023e;
    ram_cell[     198] = 32'h0;  // 32'h60fa30b2;
    ram_cell[     199] = 32'h0;  // 32'h3a81311a;
    ram_cell[     200] = 32'h0;  // 32'hf1faedaf;
    ram_cell[     201] = 32'h0;  // 32'h29b7f634;
    ram_cell[     202] = 32'h0;  // 32'h05c4fa52;
    ram_cell[     203] = 32'h0;  // 32'hc1ae9fb3;
    ram_cell[     204] = 32'h0;  // 32'ha1df77c1;
    ram_cell[     205] = 32'h0;  // 32'hb71adf3c;
    ram_cell[     206] = 32'h0;  // 32'hf1e2ecab;
    ram_cell[     207] = 32'h0;  // 32'hbd85cc0b;
    ram_cell[     208] = 32'h0;  // 32'h43e43be9;
    ram_cell[     209] = 32'h0;  // 32'h2845ba66;
    ram_cell[     210] = 32'h0;  // 32'h25cf1bb5;
    ram_cell[     211] = 32'h0;  // 32'h71cb804c;
    ram_cell[     212] = 32'h0;  // 32'h62449f05;
    ram_cell[     213] = 32'h0;  // 32'hc3f95e46;
    ram_cell[     214] = 32'h0;  // 32'h11191e16;
    ram_cell[     215] = 32'h0;  // 32'hb6b0e9b4;
    ram_cell[     216] = 32'h0;  // 32'h3b6ff463;
    ram_cell[     217] = 32'h0;  // 32'h31151ac2;
    ram_cell[     218] = 32'h0;  // 32'h2cf38072;
    ram_cell[     219] = 32'h0;  // 32'ha613f580;
    ram_cell[     220] = 32'h0;  // 32'hf72d75fe;
    ram_cell[     221] = 32'h0;  // 32'he3f771e6;
    ram_cell[     222] = 32'h0;  // 32'hd58490d7;
    ram_cell[     223] = 32'h0;  // 32'hf3fcad22;
    ram_cell[     224] = 32'h0;  // 32'h4f92c82d;
    ram_cell[     225] = 32'h0;  // 32'h38debd56;
    ram_cell[     226] = 32'h0;  // 32'h425a9edc;
    ram_cell[     227] = 32'h0;  // 32'h7b635b6a;
    ram_cell[     228] = 32'h0;  // 32'h094279c0;
    ram_cell[     229] = 32'h0;  // 32'h0729ae5f;
    ram_cell[     230] = 32'h0;  // 32'he4c8a0f5;
    ram_cell[     231] = 32'h0;  // 32'hb8ae5574;
    ram_cell[     232] = 32'h0;  // 32'h1369f03a;
    ram_cell[     233] = 32'h0;  // 32'h7dd9dcf5;
    ram_cell[     234] = 32'h0;  // 32'h7fc8be36;
    ram_cell[     235] = 32'h0;  // 32'he6322c48;
    ram_cell[     236] = 32'h0;  // 32'h1aa21641;
    ram_cell[     237] = 32'h0;  // 32'h89e06971;
    ram_cell[     238] = 32'h0;  // 32'h177db798;
    ram_cell[     239] = 32'h0;  // 32'hdff6a7e5;
    ram_cell[     240] = 32'h0;  // 32'haae5b18d;
    ram_cell[     241] = 32'h0;  // 32'h8368e85d;
    ram_cell[     242] = 32'h0;  // 32'h9370829c;
    ram_cell[     243] = 32'h0;  // 32'h4dcde27f;
    ram_cell[     244] = 32'h0;  // 32'h4c94ef3d;
    ram_cell[     245] = 32'h0;  // 32'h7fd0b2ab;
    ram_cell[     246] = 32'h0;  // 32'hc1aecff1;
    ram_cell[     247] = 32'h0;  // 32'he5947824;
    ram_cell[     248] = 32'h0;  // 32'h309180df;
    ram_cell[     249] = 32'h0;  // 32'hcd848677;
    ram_cell[     250] = 32'h0;  // 32'hce8b7bf7;
    ram_cell[     251] = 32'h0;  // 32'hee1703b5;
    ram_cell[     252] = 32'h0;  // 32'hd4e65940;
    ram_cell[     253] = 32'h0;  // 32'h84b3c6ac;
    ram_cell[     254] = 32'h0;  // 32'h4770df16;
    ram_cell[     255] = 32'h0;  // 32'he021c54b;
    // src matrix A
    ram_cell[     256] = 32'h5438ff4a;
    ram_cell[     257] = 32'h11306c47;
    ram_cell[     258] = 32'hf1ae2cf1;
    ram_cell[     259] = 32'h9c62ef0e;
    ram_cell[     260] = 32'haaac34c0;
    ram_cell[     261] = 32'h66084c75;
    ram_cell[     262] = 32'h9755ff61;
    ram_cell[     263] = 32'ha5cfadd2;
    ram_cell[     264] = 32'h31fd1bbd;
    ram_cell[     265] = 32'h8a4ae7ec;
    ram_cell[     266] = 32'hf8ba96b0;
    ram_cell[     267] = 32'hce49e621;
    ram_cell[     268] = 32'h54d589b2;
    ram_cell[     269] = 32'h6ff2aa53;
    ram_cell[     270] = 32'hf3fd513e;
    ram_cell[     271] = 32'hf37a37de;
    ram_cell[     272] = 32'hb0b5cd16;
    ram_cell[     273] = 32'h3f8f422d;
    ram_cell[     274] = 32'h89420777;
    ram_cell[     275] = 32'h0aacf044;
    ram_cell[     276] = 32'hba7c5697;
    ram_cell[     277] = 32'h7eea17c5;
    ram_cell[     278] = 32'h4f4789ed;
    ram_cell[     279] = 32'hd08bd965;
    ram_cell[     280] = 32'h7ca5a755;
    ram_cell[     281] = 32'hc5ee1079;
    ram_cell[     282] = 32'h9fe351ad;
    ram_cell[     283] = 32'h3fb15d46;
    ram_cell[     284] = 32'h962b1410;
    ram_cell[     285] = 32'h7466c8a2;
    ram_cell[     286] = 32'h1b3e5536;
    ram_cell[     287] = 32'h825cea8e;
    ram_cell[     288] = 32'h75c96243;
    ram_cell[     289] = 32'h7dce3fbf;
    ram_cell[     290] = 32'hbf78fbc4;
    ram_cell[     291] = 32'h3a643ab2;
    ram_cell[     292] = 32'h77cf8583;
    ram_cell[     293] = 32'h83689e26;
    ram_cell[     294] = 32'h16d0c224;
    ram_cell[     295] = 32'h87f400b9;
    ram_cell[     296] = 32'h3f9914bd;
    ram_cell[     297] = 32'h2d7a9ec2;
    ram_cell[     298] = 32'h7e3fcbe7;
    ram_cell[     299] = 32'h1ff8c082;
    ram_cell[     300] = 32'h625d67e0;
    ram_cell[     301] = 32'h58cbedf6;
    ram_cell[     302] = 32'hba097465;
    ram_cell[     303] = 32'h1a81f4cc;
    ram_cell[     304] = 32'hbd5dadfa;
    ram_cell[     305] = 32'h82948a08;
    ram_cell[     306] = 32'hbbde4336;
    ram_cell[     307] = 32'h086709fc;
    ram_cell[     308] = 32'hc9c9b346;
    ram_cell[     309] = 32'h1cac1db8;
    ram_cell[     310] = 32'h6efc9ca2;
    ram_cell[     311] = 32'h4f80ec4b;
    ram_cell[     312] = 32'h7e6551b4;
    ram_cell[     313] = 32'h7966e0c8;
    ram_cell[     314] = 32'hec863215;
    ram_cell[     315] = 32'hca446468;
    ram_cell[     316] = 32'hb78f5225;
    ram_cell[     317] = 32'ha7345a55;
    ram_cell[     318] = 32'ha54430c3;
    ram_cell[     319] = 32'h408f2e91;
    ram_cell[     320] = 32'h8f93ea97;
    ram_cell[     321] = 32'h83f44b49;
    ram_cell[     322] = 32'hece0481a;
    ram_cell[     323] = 32'h30dbec08;
    ram_cell[     324] = 32'ha9c6b09b;
    ram_cell[     325] = 32'h7b29d376;
    ram_cell[     326] = 32'h64639b0d;
    ram_cell[     327] = 32'h62408a4f;
    ram_cell[     328] = 32'hf6631688;
    ram_cell[     329] = 32'h5088363c;
    ram_cell[     330] = 32'h5a421e19;
    ram_cell[     331] = 32'h9a60f939;
    ram_cell[     332] = 32'hd03e934a;
    ram_cell[     333] = 32'h6f1da127;
    ram_cell[     334] = 32'hdba1094c;
    ram_cell[     335] = 32'h4327659a;
    ram_cell[     336] = 32'h13484a9a;
    ram_cell[     337] = 32'h608c00ec;
    ram_cell[     338] = 32'h214d53ec;
    ram_cell[     339] = 32'h23de7745;
    ram_cell[     340] = 32'habbf2ad0;
    ram_cell[     341] = 32'heb423178;
    ram_cell[     342] = 32'h2e83eb72;
    ram_cell[     343] = 32'hf577d9d0;
    ram_cell[     344] = 32'h6130caf3;
    ram_cell[     345] = 32'h75da0903;
    ram_cell[     346] = 32'hfedb5fe9;
    ram_cell[     347] = 32'h8c2db7a3;
    ram_cell[     348] = 32'hf1ab6a38;
    ram_cell[     349] = 32'h1645af65;
    ram_cell[     350] = 32'h0580da2c;
    ram_cell[     351] = 32'h8f0cf244;
    ram_cell[     352] = 32'h35ee647c;
    ram_cell[     353] = 32'h9e3e2754;
    ram_cell[     354] = 32'hb9f1ca9d;
    ram_cell[     355] = 32'hd69b4d78;
    ram_cell[     356] = 32'heaa19fae;
    ram_cell[     357] = 32'hd4e2de1f;
    ram_cell[     358] = 32'h804d28c4;
    ram_cell[     359] = 32'hb483b420;
    ram_cell[     360] = 32'hd7031853;
    ram_cell[     361] = 32'hd92f17d8;
    ram_cell[     362] = 32'he61e3c94;
    ram_cell[     363] = 32'h2941db36;
    ram_cell[     364] = 32'h0f4fa998;
    ram_cell[     365] = 32'h50e2cc42;
    ram_cell[     366] = 32'h290b023b;
    ram_cell[     367] = 32'h12344857;
    ram_cell[     368] = 32'h11c5208a;
    ram_cell[     369] = 32'h45b342e3;
    ram_cell[     370] = 32'h67503140;
    ram_cell[     371] = 32'hd85fdbc9;
    ram_cell[     372] = 32'h0d379d62;
    ram_cell[     373] = 32'hb025953c;
    ram_cell[     374] = 32'h694c29dd;
    ram_cell[     375] = 32'h20fe3098;
    ram_cell[     376] = 32'hc75bae82;
    ram_cell[     377] = 32'hc15cb215;
    ram_cell[     378] = 32'he8701d0b;
    ram_cell[     379] = 32'h57105f2e;
    ram_cell[     380] = 32'h25d1043e;
    ram_cell[     381] = 32'h88d9726d;
    ram_cell[     382] = 32'heac7925b;
    ram_cell[     383] = 32'hf8901f0e;
    ram_cell[     384] = 32'h468d359e;
    ram_cell[     385] = 32'h5d6d4a78;
    ram_cell[     386] = 32'h05cfef78;
    ram_cell[     387] = 32'h0e07e6b6;
    ram_cell[     388] = 32'ha1903c06;
    ram_cell[     389] = 32'hf070af66;
    ram_cell[     390] = 32'ha66a89f7;
    ram_cell[     391] = 32'h94ba4f37;
    ram_cell[     392] = 32'h28f939fd;
    ram_cell[     393] = 32'h1f885910;
    ram_cell[     394] = 32'h2b9fe4d3;
    ram_cell[     395] = 32'hac7452ad;
    ram_cell[     396] = 32'h92e18070;
    ram_cell[     397] = 32'hb793a91b;
    ram_cell[     398] = 32'h9dfc24a7;
    ram_cell[     399] = 32'h0e4d3b85;
    ram_cell[     400] = 32'habeaf7d6;
    ram_cell[     401] = 32'h6da9964c;
    ram_cell[     402] = 32'h7b026c89;
    ram_cell[     403] = 32'h381c8c64;
    ram_cell[     404] = 32'ha7e9edf8;
    ram_cell[     405] = 32'hcecf0df5;
    ram_cell[     406] = 32'h128270a0;
    ram_cell[     407] = 32'h7b1a76fc;
    ram_cell[     408] = 32'h466f8a99;
    ram_cell[     409] = 32'he1518cc1;
    ram_cell[     410] = 32'h64347ced;
    ram_cell[     411] = 32'h693d2ec9;
    ram_cell[     412] = 32'hf67899cc;
    ram_cell[     413] = 32'h10e02f9b;
    ram_cell[     414] = 32'hbdedfef5;
    ram_cell[     415] = 32'h007941b9;
    ram_cell[     416] = 32'hd5bf41aa;
    ram_cell[     417] = 32'hc96f342b;
    ram_cell[     418] = 32'hff43f741;
    ram_cell[     419] = 32'h10f3f743;
    ram_cell[     420] = 32'h6f0d05cc;
    ram_cell[     421] = 32'h3b30be5a;
    ram_cell[     422] = 32'h6c8ba858;
    ram_cell[     423] = 32'hc7c0b0d8;
    ram_cell[     424] = 32'hc98d6f3a;
    ram_cell[     425] = 32'hd32c95d7;
    ram_cell[     426] = 32'h6d947595;
    ram_cell[     427] = 32'h29492899;
    ram_cell[     428] = 32'h59d71126;
    ram_cell[     429] = 32'h900fc33c;
    ram_cell[     430] = 32'hc6271d39;
    ram_cell[     431] = 32'h5c05fbcf;
    ram_cell[     432] = 32'h6db521e5;
    ram_cell[     433] = 32'h5abab1bf;
    ram_cell[     434] = 32'hede39194;
    ram_cell[     435] = 32'h72302a57;
    ram_cell[     436] = 32'h99537906;
    ram_cell[     437] = 32'h90130219;
    ram_cell[     438] = 32'h41735542;
    ram_cell[     439] = 32'hf4f07f8c;
    ram_cell[     440] = 32'h3f85e18d;
    ram_cell[     441] = 32'hdacabbad;
    ram_cell[     442] = 32'h898f7023;
    ram_cell[     443] = 32'h3e601235;
    ram_cell[     444] = 32'h7ebd894a;
    ram_cell[     445] = 32'hd8b33aea;
    ram_cell[     446] = 32'h28b18b31;
    ram_cell[     447] = 32'hf90c756a;
    ram_cell[     448] = 32'h896bd076;
    ram_cell[     449] = 32'h2c675624;
    ram_cell[     450] = 32'h04b2492d;
    ram_cell[     451] = 32'h5d24945f;
    ram_cell[     452] = 32'ha81b0962;
    ram_cell[     453] = 32'h36b63d82;
    ram_cell[     454] = 32'hfc09641d;
    ram_cell[     455] = 32'hea9720e2;
    ram_cell[     456] = 32'hca5fe27a;
    ram_cell[     457] = 32'h644fa0d3;
    ram_cell[     458] = 32'hf3074bcf;
    ram_cell[     459] = 32'hb6113b10;
    ram_cell[     460] = 32'hc74887ba;
    ram_cell[     461] = 32'h249de0be;
    ram_cell[     462] = 32'h68f1c6ec;
    ram_cell[     463] = 32'h8823373b;
    ram_cell[     464] = 32'h784144c3;
    ram_cell[     465] = 32'h6f699c5b;
    ram_cell[     466] = 32'hdc1ec570;
    ram_cell[     467] = 32'h3e81e544;
    ram_cell[     468] = 32'hc01a21b1;
    ram_cell[     469] = 32'h27faf4bf;
    ram_cell[     470] = 32'he0909cea;
    ram_cell[     471] = 32'hfd8bca98;
    ram_cell[     472] = 32'h659990da;
    ram_cell[     473] = 32'he2dd490f;
    ram_cell[     474] = 32'hdf882114;
    ram_cell[     475] = 32'h63b452d0;
    ram_cell[     476] = 32'h2f663446;
    ram_cell[     477] = 32'haa80710a;
    ram_cell[     478] = 32'h8defc4bd;
    ram_cell[     479] = 32'hb34753fc;
    ram_cell[     480] = 32'hcbdb6200;
    ram_cell[     481] = 32'hc53b2878;
    ram_cell[     482] = 32'h0d977936;
    ram_cell[     483] = 32'hd98b910f;
    ram_cell[     484] = 32'hcf176f64;
    ram_cell[     485] = 32'h30984dae;
    ram_cell[     486] = 32'hb1325a1a;
    ram_cell[     487] = 32'h1d97469d;
    ram_cell[     488] = 32'h093de727;
    ram_cell[     489] = 32'hed598df1;
    ram_cell[     490] = 32'h69fb4c06;
    ram_cell[     491] = 32'h49afff16;
    ram_cell[     492] = 32'ha1c082d6;
    ram_cell[     493] = 32'h82dd881a;
    ram_cell[     494] = 32'h69767f97;
    ram_cell[     495] = 32'h0b704b25;
    ram_cell[     496] = 32'hd70c7b3b;
    ram_cell[     497] = 32'ha3e9e098;
    ram_cell[     498] = 32'he4c4a008;
    ram_cell[     499] = 32'h25e98b9b;
    ram_cell[     500] = 32'hd0572597;
    ram_cell[     501] = 32'h9c70053c;
    ram_cell[     502] = 32'h1df782ff;
    ram_cell[     503] = 32'h9cdc92d5;
    ram_cell[     504] = 32'h8110b82d;
    ram_cell[     505] = 32'hfaad129a;
    ram_cell[     506] = 32'hefbe8cf8;
    ram_cell[     507] = 32'h991c777a;
    ram_cell[     508] = 32'h4751a1c8;
    ram_cell[     509] = 32'ha9d45de9;
    ram_cell[     510] = 32'h93e1d87c;
    ram_cell[     511] = 32'h7c59d9f5;
    // src matrix B
    ram_cell[     512] = 32'hf6dfb51c;
    ram_cell[     513] = 32'h93d6853c;
    ram_cell[     514] = 32'hf8ef2a1c;
    ram_cell[     515] = 32'h0e9d3960;
    ram_cell[     516] = 32'h405fb9e5;
    ram_cell[     517] = 32'h6ac50477;
    ram_cell[     518] = 32'h85a5917b;
    ram_cell[     519] = 32'h51775312;
    ram_cell[     520] = 32'hb66a4ea0;
    ram_cell[     521] = 32'hb9ef24bf;
    ram_cell[     522] = 32'h03307975;
    ram_cell[     523] = 32'hea6a9012;
    ram_cell[     524] = 32'h5dd810f0;
    ram_cell[     525] = 32'h256e2311;
    ram_cell[     526] = 32'hdecd9349;
    ram_cell[     527] = 32'h301d40e5;
    ram_cell[     528] = 32'h384d43a9;
    ram_cell[     529] = 32'he7b374eb;
    ram_cell[     530] = 32'hde0d20b0;
    ram_cell[     531] = 32'h8b7c0b22;
    ram_cell[     532] = 32'h0d77aed6;
    ram_cell[     533] = 32'hf33f8ad6;
    ram_cell[     534] = 32'h763e2083;
    ram_cell[     535] = 32'h6668c126;
    ram_cell[     536] = 32'ha0f0170e;
    ram_cell[     537] = 32'hb5c0849f;
    ram_cell[     538] = 32'he74206dc;
    ram_cell[     539] = 32'h8d8c9e10;
    ram_cell[     540] = 32'h86f61de1;
    ram_cell[     541] = 32'hc17568ee;
    ram_cell[     542] = 32'h8f90aa19;
    ram_cell[     543] = 32'h66faf334;
    ram_cell[     544] = 32'h3670e364;
    ram_cell[     545] = 32'h9ff6a1f2;
    ram_cell[     546] = 32'hd18f1863;
    ram_cell[     547] = 32'h7bc31908;
    ram_cell[     548] = 32'h81c9c674;
    ram_cell[     549] = 32'h31e929f2;
    ram_cell[     550] = 32'h91226be1;
    ram_cell[     551] = 32'h1be6c771;
    ram_cell[     552] = 32'h5e5ff0dd;
    ram_cell[     553] = 32'h7ec214ae;
    ram_cell[     554] = 32'h95405d72;
    ram_cell[     555] = 32'hfbab9b51;
    ram_cell[     556] = 32'h43a37980;
    ram_cell[     557] = 32'hdaff2c35;
    ram_cell[     558] = 32'h5c1546e8;
    ram_cell[     559] = 32'ha67536d4;
    ram_cell[     560] = 32'hd6699aaa;
    ram_cell[     561] = 32'h4a3003cc;
    ram_cell[     562] = 32'h0b88205a;
    ram_cell[     563] = 32'hc9d47997;
    ram_cell[     564] = 32'h97f0af03;
    ram_cell[     565] = 32'h3770c85e;
    ram_cell[     566] = 32'h839207d5;
    ram_cell[     567] = 32'ha753dbf2;
    ram_cell[     568] = 32'h94c9b4f8;
    ram_cell[     569] = 32'h756c703e;
    ram_cell[     570] = 32'hc18222f5;
    ram_cell[     571] = 32'hdd69da77;
    ram_cell[     572] = 32'h97c11df9;
    ram_cell[     573] = 32'hc13dd686;
    ram_cell[     574] = 32'haa42d459;
    ram_cell[     575] = 32'h3988afe5;
    ram_cell[     576] = 32'hadceb040;
    ram_cell[     577] = 32'he776b97b;
    ram_cell[     578] = 32'ha78f1ac1;
    ram_cell[     579] = 32'hc0cf8bd4;
    ram_cell[     580] = 32'h47418804;
    ram_cell[     581] = 32'h4f6aea83;
    ram_cell[     582] = 32'h3555f02b;
    ram_cell[     583] = 32'h9bce053d;
    ram_cell[     584] = 32'h354deddf;
    ram_cell[     585] = 32'hd6bcec60;
    ram_cell[     586] = 32'headfa71f;
    ram_cell[     587] = 32'he37acc27;
    ram_cell[     588] = 32'h0e689f90;
    ram_cell[     589] = 32'h35342639;
    ram_cell[     590] = 32'haf55d0da;
    ram_cell[     591] = 32'h20692c88;
    ram_cell[     592] = 32'h7f846a1c;
    ram_cell[     593] = 32'h59facfeb;
    ram_cell[     594] = 32'h3fdd86a7;
    ram_cell[     595] = 32'h4007ff7c;
    ram_cell[     596] = 32'hc0955dd5;
    ram_cell[     597] = 32'hfad86ac2;
    ram_cell[     598] = 32'h3b377e07;
    ram_cell[     599] = 32'h2aa54d1f;
    ram_cell[     600] = 32'he08d47c9;
    ram_cell[     601] = 32'he154a6ed;
    ram_cell[     602] = 32'h4545d96a;
    ram_cell[     603] = 32'h6317b9dc;
    ram_cell[     604] = 32'h50bd735e;
    ram_cell[     605] = 32'hf69ab481;
    ram_cell[     606] = 32'h9fc81e02;
    ram_cell[     607] = 32'hfb2b6332;
    ram_cell[     608] = 32'h905385cb;
    ram_cell[     609] = 32'hcdef9047;
    ram_cell[     610] = 32'h8f86c538;
    ram_cell[     611] = 32'h564974e3;
    ram_cell[     612] = 32'h243b327d;
    ram_cell[     613] = 32'hb690b02f;
    ram_cell[     614] = 32'he0111218;
    ram_cell[     615] = 32'h594f7044;
    ram_cell[     616] = 32'h274c3259;
    ram_cell[     617] = 32'hb710f737;
    ram_cell[     618] = 32'hc6010bd8;
    ram_cell[     619] = 32'hb57a8fb5;
    ram_cell[     620] = 32'h6cb82b2c;
    ram_cell[     621] = 32'hdb1818c2;
    ram_cell[     622] = 32'hf19874e3;
    ram_cell[     623] = 32'h135b5b2f;
    ram_cell[     624] = 32'he7c9aded;
    ram_cell[     625] = 32'he2eb1de9;
    ram_cell[     626] = 32'hcc820784;
    ram_cell[     627] = 32'h4add16a4;
    ram_cell[     628] = 32'h79ccfd97;
    ram_cell[     629] = 32'h147c27da;
    ram_cell[     630] = 32'hfe2413bd;
    ram_cell[     631] = 32'ha105d4a8;
    ram_cell[     632] = 32'hb2ddb461;
    ram_cell[     633] = 32'h5e83309f;
    ram_cell[     634] = 32'h847a3955;
    ram_cell[     635] = 32'hdd53d9a7;
    ram_cell[     636] = 32'h015070c7;
    ram_cell[     637] = 32'ha8564dbe;
    ram_cell[     638] = 32'ha0b445f6;
    ram_cell[     639] = 32'h3140534d;
    ram_cell[     640] = 32'hcc6d3381;
    ram_cell[     641] = 32'hdb7c8c20;
    ram_cell[     642] = 32'h4f16904f;
    ram_cell[     643] = 32'hacdd2472;
    ram_cell[     644] = 32'hfc5d1599;
    ram_cell[     645] = 32'h05861c31;
    ram_cell[     646] = 32'h9b38fcb0;
    ram_cell[     647] = 32'h6eff717a;
    ram_cell[     648] = 32'h0c4af75f;
    ram_cell[     649] = 32'h9231335d;
    ram_cell[     650] = 32'h1442e79e;
    ram_cell[     651] = 32'h6a9d29ec;
    ram_cell[     652] = 32'h96d9e6f3;
    ram_cell[     653] = 32'h292b5fda;
    ram_cell[     654] = 32'h11cd49dd;
    ram_cell[     655] = 32'h2c7672ce;
    ram_cell[     656] = 32'h28e394c7;
    ram_cell[     657] = 32'h99abbc34;
    ram_cell[     658] = 32'h3da6ccaf;
    ram_cell[     659] = 32'h9d9b468c;
    ram_cell[     660] = 32'h3aa68513;
    ram_cell[     661] = 32'hc5f043c1;
    ram_cell[     662] = 32'h1854718c;
    ram_cell[     663] = 32'h45ba1f7d;
    ram_cell[     664] = 32'h6aba18cc;
    ram_cell[     665] = 32'h882f580e;
    ram_cell[     666] = 32'hffe29c3e;
    ram_cell[     667] = 32'h651928b2;
    ram_cell[     668] = 32'hc04da356;
    ram_cell[     669] = 32'hd2f20349;
    ram_cell[     670] = 32'ha4899fc3;
    ram_cell[     671] = 32'hee1ea167;
    ram_cell[     672] = 32'hdc2932f8;
    ram_cell[     673] = 32'hde7c3b80;
    ram_cell[     674] = 32'h04e012d1;
    ram_cell[     675] = 32'h2267b663;
    ram_cell[     676] = 32'h9be36598;
    ram_cell[     677] = 32'hcd031abe;
    ram_cell[     678] = 32'hc22da311;
    ram_cell[     679] = 32'hd9bf1baa;
    ram_cell[     680] = 32'hd7d0484e;
    ram_cell[     681] = 32'ha37bf051;
    ram_cell[     682] = 32'h816efa95;
    ram_cell[     683] = 32'hb404461f;
    ram_cell[     684] = 32'h241839d9;
    ram_cell[     685] = 32'he3930b18;
    ram_cell[     686] = 32'he856356f;
    ram_cell[     687] = 32'h76c82c54;
    ram_cell[     688] = 32'hd4aa1607;
    ram_cell[     689] = 32'h20e363ff;
    ram_cell[     690] = 32'he1f2a4aa;
    ram_cell[     691] = 32'h1ba9375c;
    ram_cell[     692] = 32'hbd212a30;
    ram_cell[     693] = 32'hecae60ff;
    ram_cell[     694] = 32'h4b91a4e4;
    ram_cell[     695] = 32'he8fb1033;
    ram_cell[     696] = 32'hf860595c;
    ram_cell[     697] = 32'h7ec1e417;
    ram_cell[     698] = 32'h7eda970b;
    ram_cell[     699] = 32'h4aa7cc98;
    ram_cell[     700] = 32'h8194a1ba;
    ram_cell[     701] = 32'h30aeda37;
    ram_cell[     702] = 32'hc46d77a6;
    ram_cell[     703] = 32'h8190893b;
    ram_cell[     704] = 32'h2e5397ba;
    ram_cell[     705] = 32'h7ffd4934;
    ram_cell[     706] = 32'h892030fa;
    ram_cell[     707] = 32'h6fb6487e;
    ram_cell[     708] = 32'hf536dd7e;
    ram_cell[     709] = 32'hdb076c11;
    ram_cell[     710] = 32'hffb82fa8;
    ram_cell[     711] = 32'h24b0191f;
    ram_cell[     712] = 32'hfdb5e24b;
    ram_cell[     713] = 32'h6830bc32;
    ram_cell[     714] = 32'h7b0457af;
    ram_cell[     715] = 32'h142e416a;
    ram_cell[     716] = 32'hbaee738b;
    ram_cell[     717] = 32'h68667091;
    ram_cell[     718] = 32'ha56a7b21;
    ram_cell[     719] = 32'h77863460;
    ram_cell[     720] = 32'hb6ab09d1;
    ram_cell[     721] = 32'h40ba6744;
    ram_cell[     722] = 32'h437c6162;
    ram_cell[     723] = 32'h38fdd6d8;
    ram_cell[     724] = 32'hffe5b88c;
    ram_cell[     725] = 32'hcf57b9d7;
    ram_cell[     726] = 32'h733719f8;
    ram_cell[     727] = 32'h93bb999b;
    ram_cell[     728] = 32'h89ebfe42;
    ram_cell[     729] = 32'h7870a7b9;
    ram_cell[     730] = 32'h0c51f421;
    ram_cell[     731] = 32'h1c4d47ec;
    ram_cell[     732] = 32'hfe88cfb4;
    ram_cell[     733] = 32'ha8e2d984;
    ram_cell[     734] = 32'hd4522e83;
    ram_cell[     735] = 32'had4de855;
    ram_cell[     736] = 32'h82f801ad;
    ram_cell[     737] = 32'h44872889;
    ram_cell[     738] = 32'h7b38bdc0;
    ram_cell[     739] = 32'hf09b756e;
    ram_cell[     740] = 32'hc0cbfae8;
    ram_cell[     741] = 32'h53da3da7;
    ram_cell[     742] = 32'hffbefeb4;
    ram_cell[     743] = 32'hfa464b91;
    ram_cell[     744] = 32'h84f9c74f;
    ram_cell[     745] = 32'h4e8cbf85;
    ram_cell[     746] = 32'h5a6b7586;
    ram_cell[     747] = 32'h25d05ee3;
    ram_cell[     748] = 32'hfd1b030d;
    ram_cell[     749] = 32'h628fa4ac;
    ram_cell[     750] = 32'h6fa5fd8e;
    ram_cell[     751] = 32'h3f3f4bde;
    ram_cell[     752] = 32'had0714cf;
    ram_cell[     753] = 32'hb330ff60;
    ram_cell[     754] = 32'hf4bc008a;
    ram_cell[     755] = 32'h324e01b1;
    ram_cell[     756] = 32'h58c8c944;
    ram_cell[     757] = 32'h5cc6309e;
    ram_cell[     758] = 32'h7757e33d;
    ram_cell[     759] = 32'h708320d2;
    ram_cell[     760] = 32'hf0ee87df;
    ram_cell[     761] = 32'he3c1ca64;
    ram_cell[     762] = 32'h6625f4ce;
    ram_cell[     763] = 32'h3bf146a5;
    ram_cell[     764] = 32'hfbe5cfe1;
    ram_cell[     765] = 32'hc6b628ac;
    ram_cell[     766] = 32'hca8f2fef;
    ram_cell[     767] = 32'h5a51d10a;
end

endmodule

