
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [0:768-1] [31:0] ram_cell;

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h2e23f2ec;
    ram_cell[       1] = 32'h0;  // 32'h2a25ddc0;
    ram_cell[       2] = 32'h0;  // 32'h5f810c6d;
    ram_cell[       3] = 32'h0;  // 32'hc964eeeb;
    ram_cell[       4] = 32'h0;  // 32'h6995473e;
    ram_cell[       5] = 32'h0;  // 32'hefbf23f7;
    ram_cell[       6] = 32'h0;  // 32'h69799f5f;
    ram_cell[       7] = 32'h0;  // 32'hb5c47ea5;
    ram_cell[       8] = 32'h0;  // 32'h842de83a;
    ram_cell[       9] = 32'h0;  // 32'h1e128653;
    ram_cell[      10] = 32'h0;  // 32'h14b8ced7;
    ram_cell[      11] = 32'h0;  // 32'had8718bb;
    ram_cell[      12] = 32'h0;  // 32'h1830ddec;
    ram_cell[      13] = 32'h0;  // 32'hb67fbfe0;
    ram_cell[      14] = 32'h0;  // 32'h89c1b79c;
    ram_cell[      15] = 32'h0;  // 32'h778b1991;
    ram_cell[      16] = 32'h0;  // 32'h7c155324;
    ram_cell[      17] = 32'h0;  // 32'h51af091b;
    ram_cell[      18] = 32'h0;  // 32'hfb61b46b;
    ram_cell[      19] = 32'h0;  // 32'ha70123d9;
    ram_cell[      20] = 32'h0;  // 32'hb1bc3202;
    ram_cell[      21] = 32'h0;  // 32'h8bcdd507;
    ram_cell[      22] = 32'h0;  // 32'had42bdfd;
    ram_cell[      23] = 32'h0;  // 32'h3ac6fa0d;
    ram_cell[      24] = 32'h0;  // 32'haee6e053;
    ram_cell[      25] = 32'h0;  // 32'hd0dace47;
    ram_cell[      26] = 32'h0;  // 32'h2985b53f;
    ram_cell[      27] = 32'h0;  // 32'habcd94e7;
    ram_cell[      28] = 32'h0;  // 32'h07677b7e;
    ram_cell[      29] = 32'h0;  // 32'hdc5dbb27;
    ram_cell[      30] = 32'h0;  // 32'h66b504c9;
    ram_cell[      31] = 32'h0;  // 32'h97507ec6;
    ram_cell[      32] = 32'h0;  // 32'h16161f66;
    ram_cell[      33] = 32'h0;  // 32'h21494d2f;
    ram_cell[      34] = 32'h0;  // 32'h04b157b6;
    ram_cell[      35] = 32'h0;  // 32'h837361c3;
    ram_cell[      36] = 32'h0;  // 32'h76b12f88;
    ram_cell[      37] = 32'h0;  // 32'h1bd8205e;
    ram_cell[      38] = 32'h0;  // 32'h4b6c4756;
    ram_cell[      39] = 32'h0;  // 32'h7a3593e2;
    ram_cell[      40] = 32'h0;  // 32'he34e36de;
    ram_cell[      41] = 32'h0;  // 32'hc179fe23;
    ram_cell[      42] = 32'h0;  // 32'he8ec1205;
    ram_cell[      43] = 32'h0;  // 32'h9ffd0b2a;
    ram_cell[      44] = 32'h0;  // 32'h48462c87;
    ram_cell[      45] = 32'h0;  // 32'ha95bfb88;
    ram_cell[      46] = 32'h0;  // 32'hc7a5277d;
    ram_cell[      47] = 32'h0;  // 32'h1582d187;
    ram_cell[      48] = 32'h0;  // 32'hc1a19db6;
    ram_cell[      49] = 32'h0;  // 32'h11926007;
    ram_cell[      50] = 32'h0;  // 32'h761feeb0;
    ram_cell[      51] = 32'h0;  // 32'h83644d92;
    ram_cell[      52] = 32'h0;  // 32'h54ca3e02;
    ram_cell[      53] = 32'h0;  // 32'heca8ba78;
    ram_cell[      54] = 32'h0;  // 32'h9636bf39;
    ram_cell[      55] = 32'h0;  // 32'h1fdc76e1;
    ram_cell[      56] = 32'h0;  // 32'hd6e1edfe;
    ram_cell[      57] = 32'h0;  // 32'h5ef2176d;
    ram_cell[      58] = 32'h0;  // 32'h55678137;
    ram_cell[      59] = 32'h0;  // 32'h8acea7d1;
    ram_cell[      60] = 32'h0;  // 32'hb92aa1e3;
    ram_cell[      61] = 32'h0;  // 32'hda5cfdb7;
    ram_cell[      62] = 32'h0;  // 32'h427b6ea6;
    ram_cell[      63] = 32'h0;  // 32'hcd27f5fb;
    ram_cell[      64] = 32'h0;  // 32'h5f4ea073;
    ram_cell[      65] = 32'h0;  // 32'h33fa1998;
    ram_cell[      66] = 32'h0;  // 32'h06569c76;
    ram_cell[      67] = 32'h0;  // 32'ha15883a1;
    ram_cell[      68] = 32'h0;  // 32'hfb0f7b3e;
    ram_cell[      69] = 32'h0;  // 32'hafecfcc4;
    ram_cell[      70] = 32'h0;  // 32'h0aeb40b1;
    ram_cell[      71] = 32'h0;  // 32'h8b30ec3b;
    ram_cell[      72] = 32'h0;  // 32'hf15f73fe;
    ram_cell[      73] = 32'h0;  // 32'h5efa1976;
    ram_cell[      74] = 32'h0;  // 32'haf222526;
    ram_cell[      75] = 32'h0;  // 32'h8bfebd9e;
    ram_cell[      76] = 32'h0;  // 32'h6d18eac2;
    ram_cell[      77] = 32'h0;  // 32'haf71f42b;
    ram_cell[      78] = 32'h0;  // 32'h44eb3ca6;
    ram_cell[      79] = 32'h0;  // 32'h74ab4034;
    ram_cell[      80] = 32'h0;  // 32'h1e203572;
    ram_cell[      81] = 32'h0;  // 32'h5cba4315;
    ram_cell[      82] = 32'h0;  // 32'h15efe827;
    ram_cell[      83] = 32'h0;  // 32'h85922df7;
    ram_cell[      84] = 32'h0;  // 32'h0a5c4692;
    ram_cell[      85] = 32'h0;  // 32'h16f00385;
    ram_cell[      86] = 32'h0;  // 32'h3af1636c;
    ram_cell[      87] = 32'h0;  // 32'h40faaf0c;
    ram_cell[      88] = 32'h0;  // 32'h0478e3ae;
    ram_cell[      89] = 32'h0;  // 32'h0e6ee52a;
    ram_cell[      90] = 32'h0;  // 32'h6bbd4bd3;
    ram_cell[      91] = 32'h0;  // 32'h5d91a8d1;
    ram_cell[      92] = 32'h0;  // 32'h30092469;
    ram_cell[      93] = 32'h0;  // 32'h5ada2a4f;
    ram_cell[      94] = 32'h0;  // 32'h7779a13b;
    ram_cell[      95] = 32'h0;  // 32'hcfdfda4a;
    ram_cell[      96] = 32'h0;  // 32'h3415410c;
    ram_cell[      97] = 32'h0;  // 32'hd878b860;
    ram_cell[      98] = 32'h0;  // 32'h6b8e3283;
    ram_cell[      99] = 32'h0;  // 32'hcf616f01;
    ram_cell[     100] = 32'h0;  // 32'hd1cc2580;
    ram_cell[     101] = 32'h0;  // 32'hf48e1d27;
    ram_cell[     102] = 32'h0;  // 32'hcc9dbcac;
    ram_cell[     103] = 32'h0;  // 32'h3ec91b05;
    ram_cell[     104] = 32'h0;  // 32'heccd9729;
    ram_cell[     105] = 32'h0;  // 32'ha533b71f;
    ram_cell[     106] = 32'h0;  // 32'h03eda416;
    ram_cell[     107] = 32'h0;  // 32'h3557ff33;
    ram_cell[     108] = 32'h0;  // 32'h5c8abcef;
    ram_cell[     109] = 32'h0;  // 32'hff1c2529;
    ram_cell[     110] = 32'h0;  // 32'habc0f53b;
    ram_cell[     111] = 32'h0;  // 32'h2eecf8ad;
    ram_cell[     112] = 32'h0;  // 32'hf02363a7;
    ram_cell[     113] = 32'h0;  // 32'he8f3ea91;
    ram_cell[     114] = 32'h0;  // 32'h4b4618da;
    ram_cell[     115] = 32'h0;  // 32'h6109cb4d;
    ram_cell[     116] = 32'h0;  // 32'h1288f5bf;
    ram_cell[     117] = 32'h0;  // 32'hc6943784;
    ram_cell[     118] = 32'h0;  // 32'h8382ea09;
    ram_cell[     119] = 32'h0;  // 32'h6dafde4e;
    ram_cell[     120] = 32'h0;  // 32'h8751580a;
    ram_cell[     121] = 32'h0;  // 32'h01fde381;
    ram_cell[     122] = 32'h0;  // 32'h59473152;
    ram_cell[     123] = 32'h0;  // 32'hd8ada318;
    ram_cell[     124] = 32'h0;  // 32'h28e75c97;
    ram_cell[     125] = 32'h0;  // 32'h2f0b9aa7;
    ram_cell[     126] = 32'h0;  // 32'h8ff10ac7;
    ram_cell[     127] = 32'h0;  // 32'h50c1cdb8;
    ram_cell[     128] = 32'h0;  // 32'hdd5b211b;
    ram_cell[     129] = 32'h0;  // 32'h2bb6eea1;
    ram_cell[     130] = 32'h0;  // 32'h6d5b9ce8;
    ram_cell[     131] = 32'h0;  // 32'h6087a3a0;
    ram_cell[     132] = 32'h0;  // 32'h0f7416ff;
    ram_cell[     133] = 32'h0;  // 32'h75fb2c0b;
    ram_cell[     134] = 32'h0;  // 32'h71cb1608;
    ram_cell[     135] = 32'h0;  // 32'hcc64f07c;
    ram_cell[     136] = 32'h0;  // 32'h8420dd5d;
    ram_cell[     137] = 32'h0;  // 32'hdc6ec828;
    ram_cell[     138] = 32'h0;  // 32'h219597d7;
    ram_cell[     139] = 32'h0;  // 32'h26ffc3a5;
    ram_cell[     140] = 32'h0;  // 32'h37cc8f3d;
    ram_cell[     141] = 32'h0;  // 32'h8630035a;
    ram_cell[     142] = 32'h0;  // 32'h3fc3a013;
    ram_cell[     143] = 32'h0;  // 32'hdbb58630;
    ram_cell[     144] = 32'h0;  // 32'hdde9d19f;
    ram_cell[     145] = 32'h0;  // 32'hce547647;
    ram_cell[     146] = 32'h0;  // 32'hefce9f16;
    ram_cell[     147] = 32'h0;  // 32'h721d01a9;
    ram_cell[     148] = 32'h0;  // 32'hdd26cda6;
    ram_cell[     149] = 32'h0;  // 32'hd4273120;
    ram_cell[     150] = 32'h0;  // 32'h88059666;
    ram_cell[     151] = 32'h0;  // 32'h62890cc6;
    ram_cell[     152] = 32'h0;  // 32'h891fc6d1;
    ram_cell[     153] = 32'h0;  // 32'h4e80c080;
    ram_cell[     154] = 32'h0;  // 32'hfff0d039;
    ram_cell[     155] = 32'h0;  // 32'ha7b7cb4b;
    ram_cell[     156] = 32'h0;  // 32'hd299e9f0;
    ram_cell[     157] = 32'h0;  // 32'h1f550bf6;
    ram_cell[     158] = 32'h0;  // 32'h88e9740d;
    ram_cell[     159] = 32'h0;  // 32'h7a6dafbe;
    ram_cell[     160] = 32'h0;  // 32'hc44f3c8c;
    ram_cell[     161] = 32'h0;  // 32'h5b9cd235;
    ram_cell[     162] = 32'h0;  // 32'haabef07b;
    ram_cell[     163] = 32'h0;  // 32'h9ea8d128;
    ram_cell[     164] = 32'h0;  // 32'h51167085;
    ram_cell[     165] = 32'h0;  // 32'h83fee46f;
    ram_cell[     166] = 32'h0;  // 32'h26c9027d;
    ram_cell[     167] = 32'h0;  // 32'h0283d8a2;
    ram_cell[     168] = 32'h0;  // 32'h0d4cf567;
    ram_cell[     169] = 32'h0;  // 32'hfe7dd0be;
    ram_cell[     170] = 32'h0;  // 32'ha8e8f49a;
    ram_cell[     171] = 32'h0;  // 32'hf33a533f;
    ram_cell[     172] = 32'h0;  // 32'h700c75ec;
    ram_cell[     173] = 32'h0;  // 32'h9a379ee5;
    ram_cell[     174] = 32'h0;  // 32'hacfa18b6;
    ram_cell[     175] = 32'h0;  // 32'h6b2fa4bd;
    ram_cell[     176] = 32'h0;  // 32'h1a394c81;
    ram_cell[     177] = 32'h0;  // 32'h3e502dc6;
    ram_cell[     178] = 32'h0;  // 32'h59e9604f;
    ram_cell[     179] = 32'h0;  // 32'h2d96e9e6;
    ram_cell[     180] = 32'h0;  // 32'ha98863e0;
    ram_cell[     181] = 32'h0;  // 32'h8baa6725;
    ram_cell[     182] = 32'h0;  // 32'h1cf2f50f;
    ram_cell[     183] = 32'h0;  // 32'h3e6baab3;
    ram_cell[     184] = 32'h0;  // 32'hf6708d13;
    ram_cell[     185] = 32'h0;  // 32'h00f364cc;
    ram_cell[     186] = 32'h0;  // 32'h44570cff;
    ram_cell[     187] = 32'h0;  // 32'hb3cedf06;
    ram_cell[     188] = 32'h0;  // 32'h4603af15;
    ram_cell[     189] = 32'h0;  // 32'h62ad8370;
    ram_cell[     190] = 32'h0;  // 32'hdd719064;
    ram_cell[     191] = 32'h0;  // 32'he9bd59f8;
    ram_cell[     192] = 32'h0;  // 32'h7bb940d4;
    ram_cell[     193] = 32'h0;  // 32'h728403d9;
    ram_cell[     194] = 32'h0;  // 32'ha183f0d6;
    ram_cell[     195] = 32'h0;  // 32'hc1207b88;
    ram_cell[     196] = 32'h0;  // 32'h6bdc65e6;
    ram_cell[     197] = 32'h0;  // 32'h9000398c;
    ram_cell[     198] = 32'h0;  // 32'ha5e1ba02;
    ram_cell[     199] = 32'h0;  // 32'h6cbda033;
    ram_cell[     200] = 32'h0;  // 32'h98525125;
    ram_cell[     201] = 32'h0;  // 32'h13af73ed;
    ram_cell[     202] = 32'h0;  // 32'hd5c05672;
    ram_cell[     203] = 32'h0;  // 32'h81db0099;
    ram_cell[     204] = 32'h0;  // 32'h53e3c48f;
    ram_cell[     205] = 32'h0;  // 32'hbc7a2b3f;
    ram_cell[     206] = 32'h0;  // 32'hfb2a191d;
    ram_cell[     207] = 32'h0;  // 32'h406db6b3;
    ram_cell[     208] = 32'h0;  // 32'h1ba75cf3;
    ram_cell[     209] = 32'h0;  // 32'h3f1c49a1;
    ram_cell[     210] = 32'h0;  // 32'h3e7b48d4;
    ram_cell[     211] = 32'h0;  // 32'h47ea4cd5;
    ram_cell[     212] = 32'h0;  // 32'hc4982679;
    ram_cell[     213] = 32'h0;  // 32'h23b63ec8;
    ram_cell[     214] = 32'h0;  // 32'h7426c26d;
    ram_cell[     215] = 32'h0;  // 32'h98f30c7a;
    ram_cell[     216] = 32'h0;  // 32'h51b153e6;
    ram_cell[     217] = 32'h0;  // 32'h046ed2a2;
    ram_cell[     218] = 32'h0;  // 32'h905fda0c;
    ram_cell[     219] = 32'h0;  // 32'h99a20d45;
    ram_cell[     220] = 32'h0;  // 32'hf6eb68a5;
    ram_cell[     221] = 32'h0;  // 32'h9fea1fda;
    ram_cell[     222] = 32'h0;  // 32'h7adfb382;
    ram_cell[     223] = 32'h0;  // 32'hb8db538b;
    ram_cell[     224] = 32'h0;  // 32'h5ec07e67;
    ram_cell[     225] = 32'h0;  // 32'h88e1d5ad;
    ram_cell[     226] = 32'h0;  // 32'hf83f3442;
    ram_cell[     227] = 32'h0;  // 32'hf4caf53b;
    ram_cell[     228] = 32'h0;  // 32'h0c217529;
    ram_cell[     229] = 32'h0;  // 32'h7b183119;
    ram_cell[     230] = 32'h0;  // 32'h03f888f2;
    ram_cell[     231] = 32'h0;  // 32'h92a96e89;
    ram_cell[     232] = 32'h0;  // 32'hd0e10fd4;
    ram_cell[     233] = 32'h0;  // 32'h28bbd470;
    ram_cell[     234] = 32'h0;  // 32'h8015c14a;
    ram_cell[     235] = 32'h0;  // 32'hf2403dfa;
    ram_cell[     236] = 32'h0;  // 32'h6f1bafbf;
    ram_cell[     237] = 32'h0;  // 32'hba716bd9;
    ram_cell[     238] = 32'h0;  // 32'ha314df6f;
    ram_cell[     239] = 32'h0;  // 32'h40c7fd22;
    ram_cell[     240] = 32'h0;  // 32'hed1681d8;
    ram_cell[     241] = 32'h0;  // 32'he158c970;
    ram_cell[     242] = 32'h0;  // 32'h4271f234;
    ram_cell[     243] = 32'h0;  // 32'ha95b2b67;
    ram_cell[     244] = 32'h0;  // 32'hf57372f0;
    ram_cell[     245] = 32'h0;  // 32'h1a1ff398;
    ram_cell[     246] = 32'h0;  // 32'h3c83b69e;
    ram_cell[     247] = 32'h0;  // 32'h5338c146;
    ram_cell[     248] = 32'h0;  // 32'hb8d95dfb;
    ram_cell[     249] = 32'h0;  // 32'h4ffa4e19;
    ram_cell[     250] = 32'h0;  // 32'h6c3a80a1;
    ram_cell[     251] = 32'h0;  // 32'h67d24610;
    ram_cell[     252] = 32'h0;  // 32'hc3a69297;
    ram_cell[     253] = 32'h0;  // 32'ha641dfff;
    ram_cell[     254] = 32'h0;  // 32'hc195dfd6;
    ram_cell[     255] = 32'h0;  // 32'he7e09252;
    // src matrix A
    ram_cell[     256] = 32'h0e2b2be5;
    ram_cell[     257] = 32'hb1c4d592;
    ram_cell[     258] = 32'he846b6c3;
    ram_cell[     259] = 32'ha37606d9;
    ram_cell[     260] = 32'hc0ae6b59;
    ram_cell[     261] = 32'hf697f551;
    ram_cell[     262] = 32'hf54cc58a;
    ram_cell[     263] = 32'h6a3267b3;
    ram_cell[     264] = 32'h2608f59a;
    ram_cell[     265] = 32'hd1ae19b7;
    ram_cell[     266] = 32'h72cb66ac;
    ram_cell[     267] = 32'h328e3b53;
    ram_cell[     268] = 32'h9d3f24db;
    ram_cell[     269] = 32'hc33b6254;
    ram_cell[     270] = 32'h3e01c63c;
    ram_cell[     271] = 32'hab686ca3;
    ram_cell[     272] = 32'hf8a4edd9;
    ram_cell[     273] = 32'hd313743d;
    ram_cell[     274] = 32'h9b98e08b;
    ram_cell[     275] = 32'h82bd7d1f;
    ram_cell[     276] = 32'hb20a8d0a;
    ram_cell[     277] = 32'h4e97cbee;
    ram_cell[     278] = 32'hba4bc9c8;
    ram_cell[     279] = 32'h354433e6;
    ram_cell[     280] = 32'h92304743;
    ram_cell[     281] = 32'h5b9cd399;
    ram_cell[     282] = 32'hf9101689;
    ram_cell[     283] = 32'hea4127bb;
    ram_cell[     284] = 32'h67f15301;
    ram_cell[     285] = 32'hcab29cd6;
    ram_cell[     286] = 32'h6b261ffe;
    ram_cell[     287] = 32'h84701c79;
    ram_cell[     288] = 32'h64f80517;
    ram_cell[     289] = 32'haea07c58;
    ram_cell[     290] = 32'h805c78f8;
    ram_cell[     291] = 32'h907214ec;
    ram_cell[     292] = 32'h446024f4;
    ram_cell[     293] = 32'hd92bfd5f;
    ram_cell[     294] = 32'h6d4e975a;
    ram_cell[     295] = 32'ha942a016;
    ram_cell[     296] = 32'hca2442a5;
    ram_cell[     297] = 32'ha958432c;
    ram_cell[     298] = 32'ha83bae12;
    ram_cell[     299] = 32'h75fcf394;
    ram_cell[     300] = 32'h5ec9f86a;
    ram_cell[     301] = 32'hcc085f1a;
    ram_cell[     302] = 32'h263953ae;
    ram_cell[     303] = 32'hc58fd146;
    ram_cell[     304] = 32'h7456525c;
    ram_cell[     305] = 32'hca3fd7fa;
    ram_cell[     306] = 32'h03c50247;
    ram_cell[     307] = 32'h2e015a4f;
    ram_cell[     308] = 32'h7a4c2813;
    ram_cell[     309] = 32'h0de50958;
    ram_cell[     310] = 32'hc2860ba0;
    ram_cell[     311] = 32'hdc33af3e;
    ram_cell[     312] = 32'hda6a275b;
    ram_cell[     313] = 32'h5eab137f;
    ram_cell[     314] = 32'ha2293ee9;
    ram_cell[     315] = 32'hd35d6253;
    ram_cell[     316] = 32'hb30eeef7;
    ram_cell[     317] = 32'h990db725;
    ram_cell[     318] = 32'h08d6f672;
    ram_cell[     319] = 32'h8bc83823;
    ram_cell[     320] = 32'hfd353e23;
    ram_cell[     321] = 32'hd2b10d3e;
    ram_cell[     322] = 32'hfd1aefef;
    ram_cell[     323] = 32'he239a8ae;
    ram_cell[     324] = 32'h8408df40;
    ram_cell[     325] = 32'h8e53ec48;
    ram_cell[     326] = 32'h5b256604;
    ram_cell[     327] = 32'h484103ae;
    ram_cell[     328] = 32'had82fb76;
    ram_cell[     329] = 32'he919a51a;
    ram_cell[     330] = 32'h588b061f;
    ram_cell[     331] = 32'h8a1daf2e;
    ram_cell[     332] = 32'hb96c22f9;
    ram_cell[     333] = 32'h55f2d722;
    ram_cell[     334] = 32'h0255c418;
    ram_cell[     335] = 32'h06b13e00;
    ram_cell[     336] = 32'hbaf0639d;
    ram_cell[     337] = 32'hed8e4798;
    ram_cell[     338] = 32'hae7b475a;
    ram_cell[     339] = 32'h8818ec30;
    ram_cell[     340] = 32'h44bec864;
    ram_cell[     341] = 32'h11b088a0;
    ram_cell[     342] = 32'h97e999fb;
    ram_cell[     343] = 32'h9a9176de;
    ram_cell[     344] = 32'h03e73952;
    ram_cell[     345] = 32'hc40be3fa;
    ram_cell[     346] = 32'he5d78519;
    ram_cell[     347] = 32'h58a572d4;
    ram_cell[     348] = 32'hc2b4d1d3;
    ram_cell[     349] = 32'h8ccf51cb;
    ram_cell[     350] = 32'h9a474b96;
    ram_cell[     351] = 32'h266f1ad8;
    ram_cell[     352] = 32'h01be7150;
    ram_cell[     353] = 32'h3d7663c0;
    ram_cell[     354] = 32'h7ca57bc4;
    ram_cell[     355] = 32'h3e76a51e;
    ram_cell[     356] = 32'h7cb93fcc;
    ram_cell[     357] = 32'h0a2449fe;
    ram_cell[     358] = 32'h39f63c98;
    ram_cell[     359] = 32'h57903f71;
    ram_cell[     360] = 32'h81251882;
    ram_cell[     361] = 32'hce1657fa;
    ram_cell[     362] = 32'h70da09ce;
    ram_cell[     363] = 32'h04bc5a28;
    ram_cell[     364] = 32'h1a27d283;
    ram_cell[     365] = 32'h4cd3551a;
    ram_cell[     366] = 32'h73a68cec;
    ram_cell[     367] = 32'haa399498;
    ram_cell[     368] = 32'h0188334b;
    ram_cell[     369] = 32'h6afe9144;
    ram_cell[     370] = 32'hc41b0389;
    ram_cell[     371] = 32'h82108c9d;
    ram_cell[     372] = 32'hf7151dd4;
    ram_cell[     373] = 32'h954eb9f3;
    ram_cell[     374] = 32'ha235938b;
    ram_cell[     375] = 32'h9d54dfd3;
    ram_cell[     376] = 32'hce840062;
    ram_cell[     377] = 32'hbb59d921;
    ram_cell[     378] = 32'hf4edeca0;
    ram_cell[     379] = 32'hbc28cc8c;
    ram_cell[     380] = 32'hc29e9aba;
    ram_cell[     381] = 32'hcc65f17e;
    ram_cell[     382] = 32'h72120646;
    ram_cell[     383] = 32'h468a0466;
    ram_cell[     384] = 32'hc00f81d8;
    ram_cell[     385] = 32'h3c71a107;
    ram_cell[     386] = 32'hb58936f4;
    ram_cell[     387] = 32'h33c86a3d;
    ram_cell[     388] = 32'hb0201118;
    ram_cell[     389] = 32'hf9bf7df5;
    ram_cell[     390] = 32'h359d1284;
    ram_cell[     391] = 32'h18aac16a;
    ram_cell[     392] = 32'hfb339211;
    ram_cell[     393] = 32'h49e175fd;
    ram_cell[     394] = 32'hfba462ad;
    ram_cell[     395] = 32'h8368382f;
    ram_cell[     396] = 32'haee05670;
    ram_cell[     397] = 32'h69d7ea36;
    ram_cell[     398] = 32'h17bf146a;
    ram_cell[     399] = 32'h5aebeb20;
    ram_cell[     400] = 32'h24cbab6b;
    ram_cell[     401] = 32'he2c3d442;
    ram_cell[     402] = 32'hc0e1ee88;
    ram_cell[     403] = 32'ha870b37f;
    ram_cell[     404] = 32'h3b23ed3f;
    ram_cell[     405] = 32'h10eb11a6;
    ram_cell[     406] = 32'h14d169b7;
    ram_cell[     407] = 32'hdb2a49f5;
    ram_cell[     408] = 32'hf7c845ba;
    ram_cell[     409] = 32'h8d9e0769;
    ram_cell[     410] = 32'h46b8f08a;
    ram_cell[     411] = 32'ha7eb8860;
    ram_cell[     412] = 32'hf3dc21dc;
    ram_cell[     413] = 32'h745770b6;
    ram_cell[     414] = 32'h3eb632e6;
    ram_cell[     415] = 32'h2f31082f;
    ram_cell[     416] = 32'hae287af1;
    ram_cell[     417] = 32'hea3c352c;
    ram_cell[     418] = 32'h9c5cc16d;
    ram_cell[     419] = 32'hd7bd9f62;
    ram_cell[     420] = 32'h55f34002;
    ram_cell[     421] = 32'he742f35e;
    ram_cell[     422] = 32'he987260f;
    ram_cell[     423] = 32'h5d402513;
    ram_cell[     424] = 32'h871d2860;
    ram_cell[     425] = 32'hb5f20c16;
    ram_cell[     426] = 32'h12ab1d89;
    ram_cell[     427] = 32'h4385b263;
    ram_cell[     428] = 32'hcbc6e6ab;
    ram_cell[     429] = 32'h7a1d5297;
    ram_cell[     430] = 32'hd7e2dd37;
    ram_cell[     431] = 32'hedcea9f3;
    ram_cell[     432] = 32'h9ea47c5b;
    ram_cell[     433] = 32'ha05f0474;
    ram_cell[     434] = 32'h2886d0c8;
    ram_cell[     435] = 32'ha50ec226;
    ram_cell[     436] = 32'hc1977d4b;
    ram_cell[     437] = 32'h97997cb7;
    ram_cell[     438] = 32'h8412279d;
    ram_cell[     439] = 32'h3403cc4a;
    ram_cell[     440] = 32'h209dab85;
    ram_cell[     441] = 32'h92e82d33;
    ram_cell[     442] = 32'hd60402fd;
    ram_cell[     443] = 32'h6e0d73d1;
    ram_cell[     444] = 32'hc0c19744;
    ram_cell[     445] = 32'h596e7a69;
    ram_cell[     446] = 32'h118016a2;
    ram_cell[     447] = 32'hd83597eb;
    ram_cell[     448] = 32'he30bce92;
    ram_cell[     449] = 32'h1ef76892;
    ram_cell[     450] = 32'h58673cef;
    ram_cell[     451] = 32'h7165838f;
    ram_cell[     452] = 32'haaaba93d;
    ram_cell[     453] = 32'h03b06389;
    ram_cell[     454] = 32'h1fbf08bb;
    ram_cell[     455] = 32'h85fdeb99;
    ram_cell[     456] = 32'h7c652717;
    ram_cell[     457] = 32'h2d94398f;
    ram_cell[     458] = 32'hdf70af5e;
    ram_cell[     459] = 32'h2b606960;
    ram_cell[     460] = 32'h9608e972;
    ram_cell[     461] = 32'hdb092340;
    ram_cell[     462] = 32'h71329ff0;
    ram_cell[     463] = 32'ha566907e;
    ram_cell[     464] = 32'haeab1fa5;
    ram_cell[     465] = 32'h2eecf236;
    ram_cell[     466] = 32'h6be7a414;
    ram_cell[     467] = 32'ha178f6ef;
    ram_cell[     468] = 32'hb25cda86;
    ram_cell[     469] = 32'hc2caa539;
    ram_cell[     470] = 32'h27d45ea5;
    ram_cell[     471] = 32'h48615d6c;
    ram_cell[     472] = 32'h8a40f446;
    ram_cell[     473] = 32'hecc1422c;
    ram_cell[     474] = 32'h66dc3931;
    ram_cell[     475] = 32'h75c9965f;
    ram_cell[     476] = 32'h51a11b6b;
    ram_cell[     477] = 32'h8f83b0f3;
    ram_cell[     478] = 32'h92682a11;
    ram_cell[     479] = 32'h5c4e6727;
    ram_cell[     480] = 32'h7f68b59d;
    ram_cell[     481] = 32'h150787e3;
    ram_cell[     482] = 32'h6fa587a3;
    ram_cell[     483] = 32'hbfe78692;
    ram_cell[     484] = 32'h9e48d1b7;
    ram_cell[     485] = 32'hb99c8fc5;
    ram_cell[     486] = 32'hfcd6162b;
    ram_cell[     487] = 32'h1776c5b7;
    ram_cell[     488] = 32'h38f8e0a7;
    ram_cell[     489] = 32'h52157820;
    ram_cell[     490] = 32'h74b704b1;
    ram_cell[     491] = 32'h15fa9493;
    ram_cell[     492] = 32'h9ee04466;
    ram_cell[     493] = 32'h7f606654;
    ram_cell[     494] = 32'h83ee26b8;
    ram_cell[     495] = 32'h05e2da0e;
    ram_cell[     496] = 32'hd9e513f3;
    ram_cell[     497] = 32'hb1a3e16e;
    ram_cell[     498] = 32'hb9dbfb5c;
    ram_cell[     499] = 32'h2a31493e;
    ram_cell[     500] = 32'h33d659a9;
    ram_cell[     501] = 32'h2867d4c7;
    ram_cell[     502] = 32'h8c4447a5;
    ram_cell[     503] = 32'h097a6fcd;
    ram_cell[     504] = 32'hd476312a;
    ram_cell[     505] = 32'h10691050;
    ram_cell[     506] = 32'h07851e14;
    ram_cell[     507] = 32'hc35e5c62;
    ram_cell[     508] = 32'h89a20b3e;
    ram_cell[     509] = 32'h4e239ec2;
    ram_cell[     510] = 32'h06b765fe;
    ram_cell[     511] = 32'h5218d33f;
    // src matrix B
    ram_cell[     512] = 32'h7eff4d75;
    ram_cell[     513] = 32'h0c0b3a2c;
    ram_cell[     514] = 32'h4450fe80;
    ram_cell[     515] = 32'hc24d8a22;
    ram_cell[     516] = 32'h072a8a4c;
    ram_cell[     517] = 32'ha8783d86;
    ram_cell[     518] = 32'h11a2ab75;
    ram_cell[     519] = 32'h9aeec5cf;
    ram_cell[     520] = 32'hb565649c;
    ram_cell[     521] = 32'hbc45e4cd;
    ram_cell[     522] = 32'h89f05735;
    ram_cell[     523] = 32'h528e5e6a;
    ram_cell[     524] = 32'ha4ba5766;
    ram_cell[     525] = 32'hd78b8953;
    ram_cell[     526] = 32'h80e324f6;
    ram_cell[     527] = 32'h5e69355f;
    ram_cell[     528] = 32'hf47c320f;
    ram_cell[     529] = 32'h8dbaa655;
    ram_cell[     530] = 32'h429c0716;
    ram_cell[     531] = 32'h20035c0e;
    ram_cell[     532] = 32'h8ac0d1d7;
    ram_cell[     533] = 32'h78074e37;
    ram_cell[     534] = 32'h7ffd601b;
    ram_cell[     535] = 32'h4037d8ce;
    ram_cell[     536] = 32'h7838c915;
    ram_cell[     537] = 32'hfd40f53e;
    ram_cell[     538] = 32'hd411a98d;
    ram_cell[     539] = 32'hdc7bd828;
    ram_cell[     540] = 32'h7829c7c9;
    ram_cell[     541] = 32'h7098f490;
    ram_cell[     542] = 32'h440a8623;
    ram_cell[     543] = 32'h113e8a8d;
    ram_cell[     544] = 32'h81271b07;
    ram_cell[     545] = 32'h7c9bd816;
    ram_cell[     546] = 32'hb40af2b9;
    ram_cell[     547] = 32'h55080cfd;
    ram_cell[     548] = 32'h657d4bac;
    ram_cell[     549] = 32'hed035ef1;
    ram_cell[     550] = 32'h6aecf623;
    ram_cell[     551] = 32'h92c9ad1f;
    ram_cell[     552] = 32'h0ef7e63e;
    ram_cell[     553] = 32'h2e558a10;
    ram_cell[     554] = 32'h5e0a1c06;
    ram_cell[     555] = 32'hf8a412c7;
    ram_cell[     556] = 32'h6db51894;
    ram_cell[     557] = 32'h17e36d7e;
    ram_cell[     558] = 32'h54e4ae33;
    ram_cell[     559] = 32'ha8b0246b;
    ram_cell[     560] = 32'h3a5c30f1;
    ram_cell[     561] = 32'h02da3d2f;
    ram_cell[     562] = 32'hd60cc958;
    ram_cell[     563] = 32'h93f21c9c;
    ram_cell[     564] = 32'h2fe1b8a1;
    ram_cell[     565] = 32'hbb5ef1fd;
    ram_cell[     566] = 32'hda67ee7f;
    ram_cell[     567] = 32'h81fa95a1;
    ram_cell[     568] = 32'heeeababa;
    ram_cell[     569] = 32'h66675001;
    ram_cell[     570] = 32'h03c9ad3d;
    ram_cell[     571] = 32'hffc5143a;
    ram_cell[     572] = 32'haaf598d5;
    ram_cell[     573] = 32'hd9e1953d;
    ram_cell[     574] = 32'h1dc74125;
    ram_cell[     575] = 32'h0e44b3ad;
    ram_cell[     576] = 32'hb1b683c5;
    ram_cell[     577] = 32'h520952f3;
    ram_cell[     578] = 32'he732af6e;
    ram_cell[     579] = 32'he6bfeaa6;
    ram_cell[     580] = 32'ha4350d4d;
    ram_cell[     581] = 32'hf447998d;
    ram_cell[     582] = 32'hf210baff;
    ram_cell[     583] = 32'h9ded60d7;
    ram_cell[     584] = 32'h97b94285;
    ram_cell[     585] = 32'hef50437e;
    ram_cell[     586] = 32'hf5813490;
    ram_cell[     587] = 32'had800320;
    ram_cell[     588] = 32'hef52f07b;
    ram_cell[     589] = 32'he100f165;
    ram_cell[     590] = 32'h7bd21409;
    ram_cell[     591] = 32'h4b9479c7;
    ram_cell[     592] = 32'hd8b7665c;
    ram_cell[     593] = 32'h5d4bae5e;
    ram_cell[     594] = 32'hbbb15eb2;
    ram_cell[     595] = 32'h52b44128;
    ram_cell[     596] = 32'hc39374f8;
    ram_cell[     597] = 32'h7080a767;
    ram_cell[     598] = 32'h642db7f8;
    ram_cell[     599] = 32'h40069334;
    ram_cell[     600] = 32'h01f8cada;
    ram_cell[     601] = 32'h3c56f6b5;
    ram_cell[     602] = 32'h90faea35;
    ram_cell[     603] = 32'hb24fb145;
    ram_cell[     604] = 32'hb9ca9a3c;
    ram_cell[     605] = 32'h0ef72c9d;
    ram_cell[     606] = 32'hc445d00e;
    ram_cell[     607] = 32'ha4729d31;
    ram_cell[     608] = 32'h7fd55951;
    ram_cell[     609] = 32'h33ee2331;
    ram_cell[     610] = 32'h90fc322f;
    ram_cell[     611] = 32'hcfbc97fc;
    ram_cell[     612] = 32'hb3363f02;
    ram_cell[     613] = 32'h0017aca1;
    ram_cell[     614] = 32'h228f66c3;
    ram_cell[     615] = 32'hc25637ac;
    ram_cell[     616] = 32'h1e9ff145;
    ram_cell[     617] = 32'h603fa3c1;
    ram_cell[     618] = 32'hdce2e091;
    ram_cell[     619] = 32'hbd3bfcc0;
    ram_cell[     620] = 32'h6352c978;
    ram_cell[     621] = 32'h5b62a05a;
    ram_cell[     622] = 32'h1dd3bdf7;
    ram_cell[     623] = 32'ha2263199;
    ram_cell[     624] = 32'hd866274d;
    ram_cell[     625] = 32'h99ba3175;
    ram_cell[     626] = 32'h467e7f50;
    ram_cell[     627] = 32'h379bd0c6;
    ram_cell[     628] = 32'h25e4a0db;
    ram_cell[     629] = 32'h2641fb94;
    ram_cell[     630] = 32'h3c72c4ba;
    ram_cell[     631] = 32'hbb865efc;
    ram_cell[     632] = 32'h91912cef;
    ram_cell[     633] = 32'h615c8196;
    ram_cell[     634] = 32'h5b03d4b2;
    ram_cell[     635] = 32'hbed741ec;
    ram_cell[     636] = 32'h19470384;
    ram_cell[     637] = 32'h063cfb95;
    ram_cell[     638] = 32'hac72bf40;
    ram_cell[     639] = 32'ha665d73b;
    ram_cell[     640] = 32'hf843f347;
    ram_cell[     641] = 32'ha21e4251;
    ram_cell[     642] = 32'hb513b40e;
    ram_cell[     643] = 32'h9ad0f0cb;
    ram_cell[     644] = 32'hdabff8ec;
    ram_cell[     645] = 32'h98caaf6b;
    ram_cell[     646] = 32'h25271bfb;
    ram_cell[     647] = 32'h78bcf265;
    ram_cell[     648] = 32'hd2a330bc;
    ram_cell[     649] = 32'hbec6c00f;
    ram_cell[     650] = 32'hafdfe387;
    ram_cell[     651] = 32'h5b61e66d;
    ram_cell[     652] = 32'h0c6f3fab;
    ram_cell[     653] = 32'hb1d1a0fa;
    ram_cell[     654] = 32'heb2a689b;
    ram_cell[     655] = 32'h75135351;
    ram_cell[     656] = 32'h68e23542;
    ram_cell[     657] = 32'h93d262d8;
    ram_cell[     658] = 32'h30727f68;
    ram_cell[     659] = 32'h9054c046;
    ram_cell[     660] = 32'h97944c25;
    ram_cell[     661] = 32'h7a601daa;
    ram_cell[     662] = 32'h4720a85f;
    ram_cell[     663] = 32'h7fd694d5;
    ram_cell[     664] = 32'he56c7886;
    ram_cell[     665] = 32'h95225a35;
    ram_cell[     666] = 32'hd424e6c8;
    ram_cell[     667] = 32'hf3d4e312;
    ram_cell[     668] = 32'h6d1e2664;
    ram_cell[     669] = 32'h6475c9dd;
    ram_cell[     670] = 32'hae3b369e;
    ram_cell[     671] = 32'h6fa23516;
    ram_cell[     672] = 32'h942ffc04;
    ram_cell[     673] = 32'hff2c174d;
    ram_cell[     674] = 32'h53983b38;
    ram_cell[     675] = 32'h9d6cf7cd;
    ram_cell[     676] = 32'h662f57e5;
    ram_cell[     677] = 32'h5b3dc506;
    ram_cell[     678] = 32'hb0afb6d3;
    ram_cell[     679] = 32'he0d301e6;
    ram_cell[     680] = 32'hb427803a;
    ram_cell[     681] = 32'h48556762;
    ram_cell[     682] = 32'h30188067;
    ram_cell[     683] = 32'h02224cf6;
    ram_cell[     684] = 32'hde9ba91b;
    ram_cell[     685] = 32'h2415544e;
    ram_cell[     686] = 32'h58c1145a;
    ram_cell[     687] = 32'h618cdd0e;
    ram_cell[     688] = 32'h6fac429c;
    ram_cell[     689] = 32'hba572b3d;
    ram_cell[     690] = 32'h2ce7eb2a;
    ram_cell[     691] = 32'hd8919a22;
    ram_cell[     692] = 32'h355633c1;
    ram_cell[     693] = 32'h76299ce7;
    ram_cell[     694] = 32'h28d0bafb;
    ram_cell[     695] = 32'h65051881;
    ram_cell[     696] = 32'h18f9e018;
    ram_cell[     697] = 32'h7933410e;
    ram_cell[     698] = 32'h2b81d926;
    ram_cell[     699] = 32'h02bb1a03;
    ram_cell[     700] = 32'h66cb0e7d;
    ram_cell[     701] = 32'h79b79763;
    ram_cell[     702] = 32'haf933090;
    ram_cell[     703] = 32'hbb1e36ac;
    ram_cell[     704] = 32'h840a5793;
    ram_cell[     705] = 32'haf0210b9;
    ram_cell[     706] = 32'hcb37e1e9;
    ram_cell[     707] = 32'h887f84db;
    ram_cell[     708] = 32'h3119845f;
    ram_cell[     709] = 32'h17e11fa1;
    ram_cell[     710] = 32'h2e48ef02;
    ram_cell[     711] = 32'hfe11b7df;
    ram_cell[     712] = 32'ha422f290;
    ram_cell[     713] = 32'ha3b3a22d;
    ram_cell[     714] = 32'h8717c7bc;
    ram_cell[     715] = 32'h3f557fc1;
    ram_cell[     716] = 32'h2c4ff941;
    ram_cell[     717] = 32'hf01926d4;
    ram_cell[     718] = 32'h4b31dcbf;
    ram_cell[     719] = 32'h6e8a86d4;
    ram_cell[     720] = 32'hbf76c571;
    ram_cell[     721] = 32'hd3040d7a;
    ram_cell[     722] = 32'h817ef96b;
    ram_cell[     723] = 32'h07b694d7;
    ram_cell[     724] = 32'h7daef804;
    ram_cell[     725] = 32'he1efe7df;
    ram_cell[     726] = 32'hc8d06fa3;
    ram_cell[     727] = 32'hee199abc;
    ram_cell[     728] = 32'h6b6eda29;
    ram_cell[     729] = 32'h3954fa7f;
    ram_cell[     730] = 32'h460a74fe;
    ram_cell[     731] = 32'hc8ad4934;
    ram_cell[     732] = 32'h3523c743;
    ram_cell[     733] = 32'h935e5078;
    ram_cell[     734] = 32'h6fd0ec1d;
    ram_cell[     735] = 32'hd4119fbc;
    ram_cell[     736] = 32'h9cfa7b46;
    ram_cell[     737] = 32'h7acd188b;
    ram_cell[     738] = 32'h59775572;
    ram_cell[     739] = 32'ha901915b;
    ram_cell[     740] = 32'hf250eeeb;
    ram_cell[     741] = 32'h06d25bc5;
    ram_cell[     742] = 32'h76d806ea;
    ram_cell[     743] = 32'hef6ba7da;
    ram_cell[     744] = 32'hfa6d77b2;
    ram_cell[     745] = 32'h59264ea0;
    ram_cell[     746] = 32'hf1959931;
    ram_cell[     747] = 32'h9ea3b809;
    ram_cell[     748] = 32'h90ec719e;
    ram_cell[     749] = 32'ha09da789;
    ram_cell[     750] = 32'hc22fe612;
    ram_cell[     751] = 32'h5a49ff7e;
    ram_cell[     752] = 32'h4cd71974;
    ram_cell[     753] = 32'h93313145;
    ram_cell[     754] = 32'h7aa07757;
    ram_cell[     755] = 32'h935d3351;
    ram_cell[     756] = 32'hf15cab38;
    ram_cell[     757] = 32'h3d39d7b9;
    ram_cell[     758] = 32'h3ce18a19;
    ram_cell[     759] = 32'h946a1258;
    ram_cell[     760] = 32'h0b08e542;
    ram_cell[     761] = 32'ha4495c3e;
    ram_cell[     762] = 32'h96bacf88;
    ram_cell[     763] = 32'hbb12d681;
    ram_cell[     764] = 32'h3ce84e7a;
    ram_cell[     765] = 32'h007c766d;
    ram_cell[     766] = 32'he6e33260;
    ram_cell[     767] = 32'h299a76ed;
end

endmodule

